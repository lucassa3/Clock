-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Tue Oct 10 09:49:19 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ClockFSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        IN_SW0 : IN STD_LOGIC := '0';
        IN_SW1 : IN STD_LOGIC := '0';
        FSM_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END ClockFSM;

ARCHITECTURE BEHAVIOR OF ClockFSM IS
    TYPE type_fstate IS (state0,state1,state2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_FSM_OUT : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,IN_SW0,IN_SW1,reg_FSM_OUT)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state0;
            reg_FSM_OUT <= "00";
            FSM_OUT <= "00";
        ELSE
            reg_FSM_OUT <= "00";
            FSM_OUT <= "00";
            CASE fstate IS
                WHEN state0 =>
                    IF (((IN_SW0 = '1') AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((NOT((IN_SW0 = '1')) AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state0;
                    ELSIF ((NOT((IN_SW0 = '1')) AND (IN_SW1 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;

                    reg_FSM_OUT <= "00";
                WHEN state1 =>
                    IF ((NOT((IN_SW0 = '1')) AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state0;
                    ELSIF (((IN_SW0 = '1') AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((NOT((IN_SW0 = '1')) AND (IN_SW1 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_FSM_OUT <= "01";
                WHEN state2 =>
                    IF ((NOT((IN_SW0 = '1')) AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state0;
                    ELSIF (((IN_SW0 = '1') AND NOT((IN_SW1 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((NOT((IN_SW0 = '1')) AND (IN_SW1 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    reg_FSM_OUT <= "10";
                WHEN OTHERS => 
                    reg_FSM_OUT <= "XX";
                    report "Reach undefined state";
            END CASE;
            FSM_OUT <= reg_FSM_OUT;
        END IF;
    END PROCESS;
END BEHAVIOR;
