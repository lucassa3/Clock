library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; -- use that, it's a better coding guideline


entity led is
generic(

	bits	:	integer := 8
	
	);
	
port( 

	sel			:	in std_logic;
	ula_out		:	out std_logic
	
	);

end entity;

architecture rtl of led is
begin

		ula_out <= sel;
	

end architecture;

